  Table #2              Ride        Roll        Steer       Camber L    d File 2    Camber R    d File 2    Steer L     d File 2    Steer R     d File 2  
Ride and Roll             -0.000       1.000       0.400       0.385      -0.977      -0.384       0.965     -10.868      10.844       9.966      -9.923
Ride and Roll             -0.000       1.000      -0.000      -0.427      -0.165       0.401       0.180       0.033      -0.057       0.028       0.014
Ride and Roll             -0.000       1.000      -0.400      -1.117       0.525       1.291      -0.710       9.975      -9.998     -10.877      10.920
Ride and Roll             -0.000       1.000      -0.800      -1.717       1.125       2.362      -1.781      19.476     -19.500     -23.927      23.969
Ride and Roll             -0.000       0.600      -0.800      -1.587       1.233       2.181      -1.831      19.457     -19.474     -23.951      23.975
Ride and Roll             -0.000       0.500      -0.400      -0.926       0.631       1.076      -0.784       9.952      -9.966     -10.903      10.922
Ride and Roll             -0.000       0.500      -0.000      -0.210      -0.084       0.204       0.088       0.009      -0.023       0.007       0.012
Ride and Roll             -0.000       0.500       0.400       0.623      -0.917      -0.559       0.851     -10.898      10.884       9.948      -9.929
Ride and Roll             -0.000       0.500       0.800       1.654      -1.949      -1.242       1.534     -23.937      23.923      19.444     -19.425
Ride and Roll             -0.000      -0.000       0.800       1.899      -1.899      -1.396       1.396     -23.958      23.958      19.443     -19.443
Ride and Roll             -0.000      -0.000       0.400       0.853      -0.853      -0.739       0.739     -10.910      10.910       9.943      -9.943
Ride and Roll             -0.000      -0.000      -0.000      -0.000       0.000       0.000      -0.000       0.000      -0.000       0.000       0.000
Ride and Roll             -0.000      -0.000      -0.400      -0.739       0.739       0.853      -0.853       9.943      -9.943     -10.910      10.910
Ride and Roll             -0.000      -0.000      -0.800      -1.396       1.396       1.899      -1.899      19.443     -19.443     -23.958      23.958
Ride and Roll             -0.000      -0.400      -0.800      -1.273       1.506       1.704      -1.939      19.443     -19.428     -23.943      23.931
Ride and Roll             -0.000      -0.400      -0.400      -0.594       0.828       0.669      -0.905       9.946      -9.931     -10.902      10.890
Ride and Roll             -0.000      -0.400      -0.000       0.164       0.070      -0.168      -0.068       0.004       0.011       0.006      -0.018
Ride and Roll             -0.000      -0.400       0.400       1.032      -0.798      -0.888       0.652     -10.905      10.920       9.949      -9.961
Ride and Roll             -0.000      -0.400       0.800       2.088      -1.855      -1.522       1.287     -23.958      23.973      19.450     -19.462
Ride and Roll             -0.000      -0.800       0.800       2.272      -1.807      -1.652       1.179     -23.941      23.974      19.466     -19.486
Ride and Roll             -0.000      -1.000       0.800       2.362      -1.781      -1.717       1.125     -23.927      23.969      19.476     -19.500
Ride and Roll             -0.000      -1.000       0.400       1.291      -0.710      -1.117       0.525     -10.877      10.920       9.975      -9.998
Ride and Roll             -0.000      -1.000      -0.000       0.401       0.180      -0.427      -0.165       0.028       0.014       0.033      -0.057
Ride and Roll             -0.000      -1.000      -0.400      -0.384       0.965       0.385      -0.977       9.966      -9.923     -10.868      10.844
Ride and Roll             -0.000      -1.000      -0.800      -1.093       1.674       1.401      -1.993      19.458     -19.415     -23.891      23.867
